interface dadda_if;
  logic  clk;
  logic  reset;
  logic [3:0]  A_in;
  logic [3:0]  B_in;
  logic [7:0]  p_reg_out;
endinterface
